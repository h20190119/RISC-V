module PipelineDmem(input [31:0] address, input [31:0] write_data, input read, input write ,input reset, output reg [31:0] read_data);

integer i;
  
reg [7:0] dm [60:0];

initial
begin
for(i=0; i<61; i=i+1)
begin
dm[i]=i*2; 
end
end 

always@(*)
begin
if(reset==0)
$readmemh("Data.mem",dm);
else
begin
if(write==1)
{dm[address+3],dm[address+2],dm[address+1],dm[address]}=write_data;
else if(read==1)
read_data={dm[address+3],dm[address+2],dm[address+1],dm[address]};
end
end
endmodule
